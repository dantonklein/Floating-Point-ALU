module floating_point_alu (
    input logic clk, rst,
    input logic[31:0] in1, in2, in3,
    input logic[2:0] funct3,
    input logic[6:0] funct7,
    input logic[4:0] rs2,
    output logic[31:0] out,
    output logic[2:0] exception
);


endmodule