//this is for subtraction to determine how much shifting needs to occur to normalize
module leading_zero_detection (
    input logic[26:0] sub_result,
    output logic[4:0] shift_amount
);
//typically i would parameterize this but i dont think you can parameterize a casez statement

always_comb begin
    casez(sub_result)
        27'b1??????????????????????????: shift_amount = 0;
        27'b01?????????????????????????: shift_amount = 1;
        27'b001????????????????????????: shift_amount = 2;
        27'b0001???????????????????????: shift_amount = 3;
        27'b00001??????????????????????: shift_amount = 4;
        27'b000001?????????????????????: shift_amount = 5;
        27'b0000001????????????????????: shift_amount = 6;
        27'b00000001???????????????????: shift_amount = 7;
        27'b000000001??????????????????: shift_amount = 8;
        27'b0000000001?????????????????: shift_amount = 9;
        27'b00000000001????????????????: shift_amount = 10;
        27'b000000000001???????????????: shift_amount = 11;
        27'b0000000000001??????????????: shift_amount = 12;
        27'b00000000000001?????????????: shift_amount = 13;
        27'b000000000000001????????????: shift_amount = 14;
        27'b0000000000000001???????????: shift_amount = 15;
        27'b00000000000000001??????????: shift_amount = 16;
        27'b100000000000000001?????????: shift_amount = 17;
        27'b0000000000000000001????????: shift_amount = 18;
        27'b00000000000000000001???????: shift_amount = 19;
        27'b000000000000000000001??????: shift_amount = 20;
        27'b0000000000000000000001?????: shift_amount = 21;
        27'b00000000000000000000001????: shift_amount = 22;
        27'b000000000000000000000001???: shift_amount = 23;
        27'b0000000000000000000000001??: shift_amount = 24;
        27'b00000000000000000000000001?: shift_amount = 25;
        27'b000000000000000000000000001: shift_amount = 26;
        27'b000000000000000000000000000: shift_amount = 27;
        default: shift_amount = 0;
    endcase
end

endmodule